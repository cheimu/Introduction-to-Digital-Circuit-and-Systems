// Top-level module that defines the I/Os for the DE-1 SoC board
module DE1_SoC_1 (HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, KEY, LEDR, SW);

	output logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
	output logic [9:0] LEDR;
	input logic [3:0] KEY;
	input logic [9:0] SW;
	
	// Default values, turns off the HEX displays
	assign HEX0 = 7'b1111111;
	assign HEX1 = 7'b1111111;
	assign HEX2 = 7'b1111111;
	assign HEX3 = 7'b1111111;
	assign HEX4 = 7'b1111111;
	assign HEX5 = 7'b1111111;
	
	// Logic to check if item is discounted or not,
	assign LEDR[0] = SW[8] | SW[7] & SW[9];
	// Logic to check if item is stolen or not.
	assign LEDR[1] = ~(SW[0] | SW[8] | (SW[7] & ~SW[9]));
	
endmodule