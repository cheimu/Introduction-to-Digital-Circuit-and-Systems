module clock_divider (clock, divided_clocks);
	input logic clock;
	output logic [31:0] divided_clocks;

	initial
		divided_clocks <= 0;

	always_ff @(posedge clock)
		divided_clocks <= divided_clocks + 1;
endmodule 